// `define DISPLAY_CYCLES